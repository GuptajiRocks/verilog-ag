module one(
    input A,
    output Y
);

assign Y = ~A;

endmodule