module hello;
initial 
$display("Hello Verilog");

endmodule