module one;
    intial 
        $display("Hello World");
endmodule
