module notone(
    input A,
    output Y
    );

    assign Y = ~A;

endmodule