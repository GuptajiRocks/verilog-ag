module why();
    initial 
         $display("Hello World");        
    
endmodule