module one(
    input A,
    input B,
    output Y
);

assign Y = (A || B) && (B);

endmodule